  typedef enum int {DECODE_IN = 0, DECODE_OUT = 1} decode_component_index_t;
